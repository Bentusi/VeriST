(** * CompilerState: Compiler State Management

    This module defines the state monad and utilities for the compiler.
    (To be implemented in Phase 3)
*)

Require Import STCompiler.Common.Types.
Require Import STCompiler.Syntax.AST.
Require Import STCompiler.Syntax.Bytecode.

(** Placeholder for Phase 3 implementation *)
