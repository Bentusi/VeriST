(** * Compiler: Main Compiler Implementation

    This module implements the compiler from ST AST to bytecode.
    (To be implemented in Phase 3)
*)

Require Import STCompiler.Syntax.AST.
Require Import STCompiler.Syntax.Bytecode.
Require Import STCompiler.Compiler.CompilerState.
Require Import STCompiler.Compiler.CodeGen.

(** Placeholder for Phase 3 implementation *)
