(** * SourceSemantics: Operational Semantics for ST Source Language

    This module will define the operational semantics for the
    IEC 61131-3 ST source language. (To be implemented in Phase 2)
*)

Require Import STCompiler.Common.Types.
Require Import STCompiler.Common.Values.
Require Import STCompiler.Common.Environment.
Require Import STCompiler.Syntax.AST.
Require Import STCompiler.Semantics.Operations.

(** Placeholder for Phase 2 implementation *)
